LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.utils.ALL;

PACKAGE cu_pkg IS
    CONSTANT c_CU_REGISTER_INDEX_BITS : NATURAL := 5;

    CONSTANT c_INSTRUCTION_MAX_BITS : NATURAL := 64;
    TYPE t_CU_INSTRUCTION IS (
        -- 16 bits
        NO_OP, ADD, SUB, MUL, LSHIFT, RSHIFT, TEMP1, TEMP2, TEMP3, TEMP4, MOVE,

        -- 32 bits
        LOAD, STORE, BRANCH,

        -- 48 bits
        INVALID,

        -- 64 bits
        JUMP, MOVE_I, LOAD_I
    );
    -- How many bits does the specific instruction take
    TYPE t_CU_INSTRUCTION_SIZE IS (BIT16, BIT32, BIT48, BIT64);
    CONSTANT c_CU_INSTRUCTION_SIZE_BITS : NATURAL := 2;

    CONSTANT c_CU_FIRST_16BIT_INSTRUCTION : t_CU_INSTRUCTION := NO_OP;
    CONSTANT c_CU_LAST_16BIT_INSTRUCTION : t_CU_INSTRUCTION := MOVE;
    SUBTYPE t_CU_16BIT_INSTRUCTION IS t_CU_INSTRUCTION RANGE c_CU_FIRST_16BIT_INSTRUCTION TO c_CU_LAST_16BIT_INSTRUCTION;
    CONSTANT c_CU_16BIT_INSTRUCTION_OPCODE_BITS : NATURAL := bits_required_for_vector(1 + t_CU_16BIT_INSTRUCTION'pos(c_CU_LAST_16BIT_INSTRUCTION) - t_CU_16BIT_INSTRUCTION'pos(c_CU_FIRST_16BIT_INSTRUCTION));

    CONSTANT c_CU_FIRST_32BIT_INSTRUCTION : t_CU_INSTRUCTION := LOAD;
    CONSTANT c_CU_LAST_32BIT_INSTRUCTION : t_CU_INSTRUCTION := STORE;
    SUBTYPE t_CU_32BIT_INSTRUCTION IS t_CU_INSTRUCTION RANGE c_CU_FIRST_32BIT_INSTRUCTION TO c_CU_LAST_32BIT_INSTRUCTION;
    CONSTANT c_CU_32BIT_INSTRUCTION_OPCODE_BITS : NATURAL := bits_required_for_vector(1 + t_CU_32BIT_INSTRUCTION'pos(c_CU_LAST_32BIT_INSTRUCTION) - t_CU_32BIT_INSTRUCTION'pos(c_CU_FIRST_32BIT_INSTRUCTION));

    CONSTANT c_CU_FIRST_48BIT_INSTRUCTION : t_CU_INSTRUCTION := INVALID;
    CONSTANT c_CU_LAST_48BIT_INSTRUCTION : t_CU_INSTRUCTION := INVALID;
    SUBTYPE t_CU_48BIT_INSTRUCTION IS t_CU_INSTRUCTION RANGE c_CU_FIRST_48BIT_INSTRUCTION TO c_CU_LAST_48BIT_INSTRUCTION;
    CONSTANT c_CU_48BIT_INSTRUCTION_OPCODE_BITS : NATURAL := bits_required_for_vector(1 + t_CU_48BIT_INSTRUCTION'pos(c_CU_LAST_48BIT_INSTRUCTION) - t_CU_48BIT_INSTRUCTION'pos(c_CU_FIRST_48BIT_INSTRUCTION));

    CONSTANT c_CU_FIRST_64BIT_INSTRUCTION : t_CU_INSTRUCTION := JUMP;
    CONSTANT c_CU_LAST_64BIT_INSTRUCTION : t_CU_INSTRUCTION := LOAD_I;
    SUBTYPE t_CU_64BIT_INSTRUCTION IS t_CU_INSTRUCTION RANGE c_CU_FIRST_64BIT_INSTRUCTION TO c_CU_LAST_64BIT_INSTRUCTION;
    CONSTANT c_CU_64BIT_INSTRUCTION_OPCODE_BITS : NATURAL := bits_required_for_vector(1 + t_CU_64BIT_INSTRUCTION'pos(c_CU_LAST_64BIT_INSTRUCTION) - t_CU_64BIT_INSTRUCTION'pos(c_CU_FIRST_64BIT_INSTRUCTION));

    CONSTANT c_MICRO_INSTRUCTION_COUNT : NATURAL := 32;
    TYPE t_CU_MICRO_INSTRUCTION IS (
        RAM_ADDRESS_IN, RAM_ADDRESS_OUT, RAM_DATA_IN, RAM_DATA_OUT,
        REGISTER_INSTRUCTION_IN, REGISTER_INSTRUCTION_OUT,
        ALU_OUT, ALU_SUBTRACT, ALU_MULTIPLY,

        --REGISTER_DATA_BUS_TO_ADDRESS_BUS_IN, REGISTER_DATA_BUS_TO_ADDRESS_BUS_OUT, REGISTER_ADDRESS_BUS_ADDER_IN, REGISTER_ADDRESS_BUS_ADDER_OUT,

        --GP_REGISTER_CONNECTED_TO_ALU_IN, GENERAL_PURPOSE_REGISTER_3_IN,
        --GP_REGISTER_CONNECTED_TO_ALU_OUT, GENERAL_PURPOSE_REGISTER_3_OUT,

        GP_REGISTER_TO_WRITE_IN, GP_REGISTER_CONNECTED_TO_DATA_BUS_OUT,
        IMMEDIATE_VALUE_CONNECTED_TO_DATA_BUS_OUT,

        PROGRAM_COUNTER_IN, PROGRAM_COUNTER_OUT, PROGRAM_COUNTER_ADDED_IN);

    CONSTANT c_MAX_MICRO_INSTRUCTION_COUNT_IN_INSTRUCTION : NATURAL := 5;

    FUNCTION get_instruction_size(signal_vector : STD_LOGIC_VECTOR) RETURN t_CU_INSTRUCTION_SIZE;
    FUNCTION to_CU_INSTRUCTION(signal_vector : STD_LOGIC_VECTOR) RETURN t_CU_INSTRUCTION;
    FUNCTION from_CU_INSTRUCTION(instruction : t_CU_INSTRUCTION) RETURN STD_LOGIC_VECTOR;
    FUNCTION convert(micro_operation : t_CU_MICRO_INSTRUCTION) RETURN STD_LOGIC_VECTOR;
END PACKAGE cu_pkg;

PACKAGE BODY cu_pkg IS
    FUNCTION get_instruction_size(signal_vector : STD_LOGIC_VECTOR) RETURN t_CU_INSTRUCTION_SIZE IS
    BEGIN
        RETURN t_CU_INSTRUCTION_SIZE'VAL(to_integer(unsigned(signal_vector(c_CU_INSTRUCTION_SIZE_BITS - 1 DOWNTO 0))));
    END FUNCTION;

    FUNCTION to_CU_INSTRUCTION(signal_vector : STD_LOGIC_VECTOR) RETURN t_CU_INSTRUCTION IS
    BEGIN
        CASE get_instruction_size(signal_vector) IS
            WHEN BIT16 => RETURN t_CU_16BIT_INSTRUCTION'VAL(to_integer(unsigned(signal_vector(c_CU_16BIT_INSTRUCTION_OPCODE_BITS + c_CU_INSTRUCTION_SIZE_BITS - 1 DOWNTO c_CU_INSTRUCTION_SIZE_BITS))));
            WHEN BIT32 => RETURN t_CU_32BIT_INSTRUCTION'VAL(t_CU_32BIT_INSTRUCTION'POS(c_CU_FIRST_32BIT_INSTRUCTION) + to_integer(unsigned(signal_vector(c_CU_32BIT_INSTRUCTION_OPCODE_BITS + c_CU_INSTRUCTION_SIZE_BITS - 1 DOWNTO c_CU_INSTRUCTION_SIZE_BITS))));
            WHEN BIT48 => RETURN t_CU_48BIT_INSTRUCTION'VAL(t_CU_48BIT_INSTRUCTION'POS(c_CU_FIRST_48BIT_INSTRUCTION) + to_integer(unsigned(signal_vector(c_CU_48BIT_INSTRUCTION_OPCODE_BITS + c_CU_INSTRUCTION_SIZE_BITS - 1 DOWNTO c_CU_INSTRUCTION_SIZE_BITS))));
            WHEN BIT64 => RETURN t_CU_64BIT_INSTRUCTION'VAL(t_CU_64BIT_INSTRUCTION'POS(c_CU_FIRST_64BIT_INSTRUCTION) + to_integer(unsigned(signal_vector(c_CU_64BIT_INSTRUCTION_OPCODE_BITS + c_CU_INSTRUCTION_SIZE_BITS - 1 DOWNTO c_CU_INSTRUCTION_SIZE_BITS))));
        END CASE;
    END FUNCTION;

    FUNCTION from_CU_INSTRUCTION(instruction : t_CU_INSTRUCTION) RETURN STD_LOGIC_VECTOR IS
    BEGIN
        IF instruction >= c_CU_FIRST_16BIT_INSTRUCTION AND instruction <= c_CU_LAST_16BIT_INSTRUCTION THEN
            RETURN (STD_LOGIC_VECTOR(to_unsigned(t_CU_16BIT_INSTRUCTION'POS(instruction), c_CU_16BIT_INSTRUCTION_OPCODE_BITS)) & STD_LOGIC_VECTOR(to_unsigned(t_CU_INSTRUCTION_SIZE'POS(BIT16), 2)));
            ELSIF instruction >= c_CU_FIRST_32BIT_INSTRUCTION AND instruction <= c_CU_LAST_32BIT_INSTRUCTION THEN
            RETURN (STD_LOGIC_VECTOR(to_unsigned(t_CU_32BIT_INSTRUCTION'POS(instruction) - t_CU_32BIT_INSTRUCTION'POS(c_CU_FIRST_32BIT_INSTRUCTION), c_CU_32BIT_INSTRUCTION_OPCODE_BITS)) & STD_LOGIC_VECTOR(to_unsigned(t_CU_INSTRUCTION_SIZE'POS(BIT32), 2)));
            ELSIF instruction >= c_CU_FIRST_48BIT_INSTRUCTION AND instruction <= c_CU_LAST_48BIT_INSTRUCTION THEN
            RETURN (STD_LOGIC_VECTOR(to_unsigned(t_CU_48BIT_INSTRUCTION'POS(instruction) - t_CU_48BIT_INSTRUCTION'POS(c_CU_FIRST_48BIT_INSTRUCTION), c_CU_48BIT_INSTRUCTION_OPCODE_BITS)) & STD_LOGIC_VECTOR(to_unsigned(t_CU_INSTRUCTION_SIZE'POS(BIT48), 2)));
            ELSE
            RETURN (STD_LOGIC_VECTOR(to_unsigned(t_CU_64BIT_INSTRUCTION'POS(instruction) - t_CU_64BIT_INSTRUCTION'POS(c_CU_FIRST_64BIT_INSTRUCTION), c_CU_64BIT_INSTRUCTION_OPCODE_BITS)) & STD_LOGIC_VECTOR(to_unsigned(t_CU_INSTRUCTION_SIZE'POS(BIT64), 2)));
        END IF;
    END FUNCTION;

    FUNCTION convert(micro_operation : t_CU_MICRO_INSTRUCTION) RETURN STD_LOGIC_VECTOR IS
    BEGIN
        RETURN STD_LOGIC_VECTOR(to_unsigned(2 ** t_CU_MICRO_INSTRUCTION'POS(micro_operation), c_MICRO_INSTRUCTION_COUNT));
    END FUNCTION;
END PACKAGE BODY cu_pkg;